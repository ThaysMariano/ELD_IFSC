-- biblioteca

package moecke is

	type integer_vector is array(natural range <>) of integer range 0 to 31;

end package;
